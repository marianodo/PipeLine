`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:47:18 01/20/2015 
// Design Name: 
// Module Name:    ControlUnit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ControlUnit(
	input [5:0] inOpcode, inFunction, //Opcode y Funcion
	input clk,
	output reg RegDst,Branch,MemRead,MemtoReg,MemWrite,ALUSrc,RegWrite,flagBranch,
	output reg [1:0] ALUOp,
	output reg [2:0] flagLoadWordDividerMEM,
	output reg [1:0] flagStoreWordDividerMEM,
	output reg [5:0] outFunction
    );
	 reg opCode;
	 
initial
begin
	RegDst = 1; // Mux para elegir Rd o Rt, en 1 elige Rd
	Branch = 0; // Es el and con el Zero de la alu
	MemtoReg = 0; //Mux que elige entre Alu o Memoria, 0 es ALU
	MemRead = 0; //Flag para leer en memoria, en 0 no pasa nada, en 1 Lee
	MemWrite = 0; //Flag para escribir en memoria, en 0 no pasa nada, en 1 Escribe
	ALUSrc = 0; //Mux que elige entre Inmediato o Rt, 1 es inmediato, 0 Rt
	RegWrite = 0; //Flag que lee o escribe en registros , 0 Lee 1 Escribe
	ALUOp = 2'b10;
	flagLoadWordDividerMEM = 0;
	flagStoreWordDividerMEM = 0;
	flagBranch = 0; // 0 = BNE, 1 = BEQ
end

always @(*)
begin
	if(clk)
		begin
			if ( inOpcode == 0) //Write R-Type
				begin
					RegDst = 1;
					Branch = 0;
					MemtoReg = 0;
					MemRead = 0;
					MemWrite = 0;
					ALUSrc = 0;
					RegWrite = 1;
					ALUOp = 2'b10;
					flagLoadWordDividerMEM = 0;
					flagStoreWordDividerMEM = 0;
					outFunction = inFunction; //Si es tipo R la funcion es igual a la funcion
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
			else if (inOpcode == 35 ) //Write Load, LW
				begin
					RegDst = 0;
					Branch = 0;
					MemtoReg = 1;
					MemRead = 0;
					MemWrite = 0;
					ALUSrc = 1;
					RegWrite = 1;
					ALUOp = 2'b00;
					flagLoadWordDividerMEM = 0;
					flagStoreWordDividerMEM = 0;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
			else if (inOpcode == 39 ) //Write Load, LWU
				begin
					RegDst = 0;
					Branch = 0;
					MemtoReg = 1;
					MemRead = 0;
					MemWrite = 0;
					ALUSrc = 1;
					RegWrite = 1;
					ALUOp = 2'b00;
					flagLoadWordDividerMEM = 1;
					flagStoreWordDividerMEM = 0;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
			else if (inOpcode == 32 ) //Write Load, LB
				begin
					RegDst = 0;
					Branch = 0;
					MemtoReg = 1;
					MemRead = 0;
					MemWrite = 0;
					ALUSrc = 1;
					RegWrite = 1;
					ALUOp = 2'b00;
					flagLoadWordDividerMEM = 2;
					flagStoreWordDividerMEM = 0;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
			else if (inOpcode == 36 ) //Write Load, LBU
				begin
					RegDst = 0;
					Branch = 0;
					MemtoReg = 1;
					MemRead = 0;
					MemWrite = 0;
					ALUSrc = 1;
					RegWrite = 1;
					ALUOp = 2'b00;
					flagLoadWordDividerMEM = 3;
					flagStoreWordDividerMEM = 0;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
			else if (inOpcode == 33 ) //Write Load, LH
				begin
					RegDst = 0;
					Branch = 0;
					MemtoReg = 1;
					MemRead = 0;
					MemWrite = 0;
					ALUSrc = 1;
					RegWrite = 1;
					ALUOp = 2'b00;
					flagLoadWordDividerMEM = 4;
					flagStoreWordDividerMEM = 0;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
			else if (inOpcode == 37 ) //Write Load, LHU
				begin
					RegDst = 0;
					Branch = 0;
					MemtoReg = 1;
					MemRead = 0;
					MemWrite = 0;
					ALUSrc = 1;
					RegWrite = 1;
					ALUOp = 2'b00;
					flagLoadWordDividerMEM = 5;
					flagStoreWordDividerMEM = 0;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
			else if (inOpcode == 43 ) //Write Store, SW
				begin
					RegDst = 0;
					Branch = 0;
					MemtoReg = 0;
					MemRead = 0;
					MemWrite = 1;
					ALUSrc = 1;
					RegWrite = 0;
					ALUOp = 2'b00;
					flagLoadWordDividerMEM = 0;
					flagStoreWordDividerMEM = 0;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
			else if (inOpcode == 40 ) //Write Store, SB
				begin
					RegDst = 0;
					Branch = 0;
					MemtoReg = 0;
					MemRead = 0;
					MemWrite = 1;
					ALUSrc = 1;
					RegWrite = 0;
					ALUOp = 2'b00;
					flagLoadWordDividerMEM = 0;
					flagStoreWordDividerMEM = 1;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
			else if (inOpcode == 41 ) //Write Store, SH
				begin
					RegDst = 0;
					Branch = 0;
					MemtoReg = 0;
					MemRead = 0;
					MemWrite = 1;
					ALUSrc = 1;
					RegWrite = 0;
					ALUOp = 2'b00;
					flagLoadWordDividerMEM = 0;
					flagStoreWordDividerMEM = 2;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
			else if (inOpcode == 4 ) //Write Branch, BEQ
				begin
					RegDst = 0;
					Branch = 1;
					MemtoReg = 0;
					MemRead = 0;
					MemWrite = 0;
					ALUSrc = 0;
					RegWrite = 0;
					ALUOp = 2'b01;
					flagLoadWordDividerMEM = 0;
					flagStoreWordDividerMEM = 0;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 1; // 0 = BNE, 1 = BEQ
				end
			else if (inOpcode == 5 ) //Write Branch, BNE
				begin
					RegDst = 0;
					Branch = 1;
					MemtoReg = 0;
					MemRead = 0;
					MemWrite = 0;
					ALUSrc = 0;
					RegWrite = 0;
					ALUOp = 2'b01;
					flagLoadWordDividerMEM = 0;
					flagStoreWordDividerMEM = 0;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
			else //El resto son inmediatas
				begin
					RegDst = 0;
					Branch = 0;
					MemtoReg = 0;
					MemRead = 0;
					MemWrite = 0;
					ALUSrc = 1;
					RegWrite = 1;
					ALUOp = 2'b11;
					flagLoadWordDividerMEM = 0;
					flagStoreWordDividerMEM = 0;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
		end
	else if(clk == 0)//Clock en 0
		begin
			if ( inOpcode == 0) //Read R-Type
				begin
					RegDst = 1;
					Branch = 0;
					MemtoReg = 0;
					MemRead = 0;
					MemWrite = 0;
					ALUSrc = 0;
					RegWrite = 0;
					ALUOp = 2'b10;
					flagLoadWordDividerMEM = 0;
					flagStoreWordDividerMEM = 0;
					outFunction = inFunction; 
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
			else if (inOpcode == 35 ) //Read Load, LW
				begin
					RegDst = 0;
					Branch = 0;
					MemtoReg = 1;
					MemRead = 1;
					MemWrite = 0;
					ALUSrc = 1;
					RegWrite = 0;
					ALUOp = 2'b00;
					flagLoadWordDividerMEM = 0;
					flagStoreWordDividerMEM = 0;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
			else if (inOpcode == 39 ) //Read Load, LWU
				begin
					RegDst = 0;
					Branch = 0;
					MemtoReg = 1;
					MemRead = 1;
					MemWrite = 0;
					ALUSrc = 1;
					RegWrite = 0;
					ALUOp = 2'b00;
					flagLoadWordDividerMEM = 1;
					flagStoreWordDividerMEM = 0;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
			else if (inOpcode == 32 ) //Read Load, LB
				begin
					RegDst = 0;
					Branch = 0;
					MemtoReg = 1;
					MemRead = 1;
					MemWrite = 0;
					ALUSrc = 1;
					RegWrite = 0;
					ALUOp = 2'b00;
					flagLoadWordDividerMEM = 2;
					flagStoreWordDividerMEM = 0;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
			else if (inOpcode == 36 ) //Read Load, LBU
				begin
					RegDst = 0;
					Branch = 0;
					MemtoReg = 1;
					MemRead = 1;
					MemWrite = 0;
					ALUSrc = 1;
					RegWrite = 0;
					ALUOp = 2'b00;
					flagLoadWordDividerMEM = 3;
					flagStoreWordDividerMEM = 0;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
			else if (inOpcode == 33 ) //Read Load, LH
				begin
					RegDst = 0;
					Branch = 0;
					MemtoReg = 1;
					MemRead = 1;
					MemWrite = 0;
					ALUSrc = 1;
					RegWrite = 0;
					ALUOp = 2'b00;
					flagLoadWordDividerMEM = 4;
					flagStoreWordDividerMEM = 0;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
			else if (inOpcode == 37 ) //Read Load, LHU
				begin
					RegDst = 0;
					Branch = 0;
					MemtoReg = 1;
					MemRead = 1;
					MemWrite = 0;
					ALUSrc = 1;
					RegWrite = 0;
					ALUOp = 2'b00;
					flagLoadWordDividerMEM = 5;
					flagStoreWordDividerMEM = 0;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
			else if (inOpcode == 43 ) //Read Store, SW
				begin
					RegDst = 0;
					Branch = 0;
					MemtoReg = 0;
					MemRead = 0;
					MemWrite = 0;
					ALUSrc = 1;
					RegWrite = 0;
					ALUOp = 2'b00;
					flagLoadWordDividerMEM = 0;
					flagStoreWordDividerMEM = 0;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
			else if (inOpcode == 40 ) //Read Store, SB
				begin
					RegDst = 0;
					Branch = 0;
					MemtoReg = 0;
					MemRead = 0;
					MemWrite = 0;
					ALUSrc = 1;
					RegWrite = 0;
					ALUOp = 2'b00;
					flagLoadWordDividerMEM = 0;
					flagStoreWordDividerMEM = 1;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
			else if (inOpcode == 41 ) //Read Store, SH
				begin
					RegDst = 1;
					Branch = 0;
					MemtoReg = 0;
					MemRead = 0;
					MemWrite = 0;
					ALUSrc = 1;
					RegWrite = 0;
					ALUOp = 2'b00;
					flagLoadWordDividerMEM = 0;
					flagStoreWordDividerMEM = 2;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
			else if (inOpcode == 4 ) //Branch, BEQ
				begin
					RegDst = 0;
					Branch = 1;
					MemtoReg = 0;
					MemRead = 0;
					MemWrite = 0;
					ALUSrc = 0;
					RegWrite = 0;
					ALUOp = 2'b01;
					flagLoadWordDividerMEM = 0;
					flagStoreWordDividerMEM = 0;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 1; // 0 = BNE, 1 = BEQ
				end
			else if (inOpcode == 5 ) //Branch, BNE
				begin
					RegDst = 0;
					Branch = 1;
					MemtoReg = 0;
					MemRead = 0;
					MemWrite = 0;
					ALUSrc = 0;
					RegWrite = 0;
					ALUOp = 2'b01;
					flagLoadWordDividerMEM = 0;
					flagStoreWordDividerMEM = 0;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
			
			else //El resto son inmediatas
				begin
					RegDst = 0;
					Branch = 0;
					MemtoReg = 0;
					MemRead = 0;
					MemWrite = 0;
					ALUSrc = 1;
					RegWrite = 0;
					ALUOp = 2'b10;
					flagLoadWordDividerMEM = 0;
					flagStoreWordDividerMEM = 0;
					outFunction = inOpcode; // Si no es r-Type, la funcion es igual al opcode
					flagBranch = 0; // 0 = BNE, 1 = BEQ
				end
		
		end
	
end

endmodule

