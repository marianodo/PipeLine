`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:32:44 01/20/2015 
// Design Name: 
// Module Name:    StageIF 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module StageIF(
    );
	 
	 
//wire [4:0] rs;
//wire [4:0] rd;
//wire [4:0] rt;
//wire [4:0] sa;
//wire [5:0] instReg;
//wire [31:0] writeData;
////wire wdSelect;
////wire [31:0] dataRd, dataRt;
//reg select = 0; 
//
//	muxPc callMuxPc (
//	.inMuxAddPc(PostPc),
//	.inMuxAddJmp(jmpAddr),
//	.select(btnSelect),
//	.outMuxPc(PcMux)
//	);
//
//	Pc callPc (
//	.inPc(PcMux),
//	.outPc(Pc)
//	);
//
//	addPc callAddPc (
//	.btn(btn),
//	.inAddPc(Pc),
//	.outAddPc(PostPc)
//	);
//	
//	InstructionMem callInstruccionMem (
//	.inInstructionMem(Pc),
//	.rsReg(rs),
//	.rtReg(rt),
//	.rdReg(rd),
//	.saReg(sa),
//	.instRreg(instReg)
//	);
	


endmodule
